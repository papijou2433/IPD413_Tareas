** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/IHP/MOS_testing/DC_hv_nmos.sch
**.subckt DC_hv_nmos vg vd vd
*.ipin vg
*.ipin vd
*.ipin vd
XM1 vd vg GND GND sg13_hv_nmos w=1.0u l=0.45u ng=1 m=1
XM2 GND vg vd vd sg13_hv_pmos w=1.0u l=0.45u ng=1 m=1
**** begin user architecture code


vgs vg 0 3.3
vds vd 0 3.3
.control
save all
save @n.xm1.nsg13_hv_nmos[ids]
save @n.xm1.nsg13_hv_nmos[vth]
save @n.xm2.nsg13_hv_pmos[ids]
save @n.xm2.nsg13_hv_pmos[vth]

dc vgs 0.0 3.3 0.05
let idn  = @n.xm1.nsg13_hv_nmos[ids]
let vthn = @n.xm1.nsg13_hv_nmos[vth]
let idp  = @n.xm2.nsg13_hv_pmos[ids]
let vthp = @n.xm2.nsg13_hv_pmos[vth]

print vthn vthp
plot idn
plot -idp

.endc


 .lib cornerMOShv.lib mos_tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
