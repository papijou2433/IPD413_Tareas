** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/IPD413_202501/xschem/Tareas/Tarea_1/cs_amp_full_IPD413HW1.sch
**.subckt cs_amp_full_IPD413HW1 vg vout
*.iopin vg
*.iopin vout
I1 VDD vout {Ids}
XM1 vout vg GND GND sg13_lv_nmos w={W} l={L} ng=1 m={mult}
**** begin user architecture code


.param corner=0

.if (corner==0)
.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ
.endif



.option wnflag=1
.param gm    = {3.1415*1.1m}
.param gm_id = 13
.param Ids   = {gm/gm_id}
.param L     = 0.13u
.param W     = 3.13u
.param mult  = 10

vsup VDD 0 1.8
vin vg 0 dc=0.45 ac=1

cload vout 0 5p

.control
save all
op
save @n.xm1.nsg13_lv_nmos[gm]
save @n.xm1.nsg13_lv_nmos[ids]
save @n.xm1.nsg13_lv_nmos[gds]
save @n.xm1.nsg13_lv_nmos[ib]

*dc vin -0.01 0.01 0.001
dc vin 0.45 0.45 0.001

let gdsn = @n.xm1.nsg13_lv_nmos[gds]
let gmn = @n.xm1.nsg13_lv_nmos[gm]
let vthn = @n.xm1.nsg13_lv_nmos[vth]
let idn = @n.xm1.nsg13_lv_nmos[ids]
let ao = gmn / gdsn

print Ao

ac dec 100 1 1T
plot vdb(vout)
meas ac GBW when vdb(vout)=0
meas ac DCG find vdb(vout) at=1]]
wrdata cs_amp_bode.raw vdb(vout)
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
